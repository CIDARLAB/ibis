/*
 And gate
*/
module and_gate
(
 input a,
 input b,
 output out
 );

   assign out = a & b;

endmodule // and_gate
